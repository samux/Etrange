module fifo (
	wire data_in[31:0],
	wire w_e,
	reg data_out[31:0],
	wire r_e);






endmodule;
